interface interf (input wclk,rclk,wreset,rreset,we,re);
logic [7:0] datain;
logic  full,empty;
logic [7:0] dataout;
endinterface
