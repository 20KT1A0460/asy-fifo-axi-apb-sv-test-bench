interface interf (input clk,reset);
logic wr;
logic [9:0] addr;
logic [15:0] datain;
logic [15:0] dataout;
endinterface
