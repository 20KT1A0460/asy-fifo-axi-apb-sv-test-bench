module endmodule
